//Copyright (C)2014-2021 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8
//Part Number: GW1NR-LV9QN88C6/I5
//Device: GW1NR-9
//Created Time: Sun Jan  9 21:01:54 2022

module Gowin_pROM (dout, clk, oce, ce, reset, ad);

output [127:0] dout;
input clk;
input oce;
input ce;
input reset;
input [6:0] ad;

wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO(dout[31:0]),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({gw_gnd,gw_gnd,ad[6:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 32;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h0000000018000000180000000000000000000000FF7E0000817E000000000000;
defparam prom_inst_0.INIT_RAM_01 = 256'h18000000637F0000333F0000663C00000E1E0000FFFFFFFF00000000FFFFFFFF;
defparam prom_inst_0.INIT_RAM_02 = 256'h3C1800000000000060C67C00DB7F0000666600003C1800000E060200E0C08000;
defparam prom_inst_0.INIT_RAM_03 = 256'h000000000000000000000000000000000000000000000000181800003C180000;
defparam prom_inst_0.INIT_RAM_04 = 256'h303030006C38000000000000C67C18186C000000666666003C18000000000000;
defparam prom_inst_0.INIT_RAM_05 = 256'h00000000000000000000000000000000000000000000000018300000180C0000;
defparam prom_inst_0.INIT_RAM_06 = 256'hC6FE000060380000C0FE00001C0C0000C67C0000C67C000038180000C67C0000;
defparam prom_inst_0.INIT_RAM_07 = 256'hC67C00006000000000000000060000000000000000000000C67C0000C67C0000;
defparam prom_inst_0.INIT_RAM_08 = 256'h663C000066FE000066FE00006CF80000663C000066FC000038100000C67C0000;
defparam prom_inst_0.INIT_RAM_09 = 256'hC67C0000E6C60000E7C3000060F0000066E600000C1E0000183C0000C6C60000;
defparam prom_inst_0.INIT_RAM_0A = 256'hC3C30000C3C30000C6C60000DBFF0000C67C000066FC0000C67C000066FC0000;
defparam prom_inst_0.INIT_RAM_0B = 256'h00000000C66C38100C3C000080000000303C0000C3FF0000C3C30000C3C30000;
defparam prom_inst_0.INIT_RAM_0C = 256'h000000006C380000000000000C1C00000000000060E000000000000000183030;
defparam prom_inst_0.INIT_RAM_0D = 256'h0000000000000000000000001838000060E00000060600001818000060E00000;
defparam prom_inst_0.INIT_RAM_0E = 256'h0000000000000000000000003010000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0F = 256'h00000000DC7600001870000018180000180E0000000000000000000000000000;

pROM prom_inst_1 (
    .DO(dout[63:32]),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({gw_gnd,gw_gnd,ad[6:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 32;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'h3C180000FFFF7E3CE7E73C3CFE7C3810FEFEFE6CC3FFFFDBBD8181A500000000;
defparam prom_inst_1.INIT_RAM_01 = 256'hE73CDB186363637F3030303F3C666666CC78321ABD99C3FF42663C00C3E7FFFF;
defparam prom_inst_1.INIT_RAM_02 = 256'h1818187E00000000C6C66C381B7BDBDB666666661818187E3EFE3E1EF8FEF8F0;
defparam prom_inst_1.INIT_RAM_03 = 256'h7C7CFEFE7C383810FF662400C0C00000FE603000FE0C1800181818181818187E;
defparam prom_inst_1.INIT_RAM_04 = 256'h00000060DC76386C180CC6C2067CC0C26C6CFE6C0000002418183C3C00000000;
defparam prom_inst_1.INIT_RAM_05 = 256'h180C0602000000007E000000000000007E181800FF3C66000C0C0C0C30303030;
defparam prom_inst_1.INIT_RAM_06 = 256'h180C0606C6FCC0C006FCC0C0FECC6C3C063C060630180C0618181878F6DECEC6;
defparam prom_inst_1.INIT_RAM_07 = 256'h18180CC6060C183000007E006030180C0000181800001818067EC6C6C67CC6C6;
defparam prom_inst_1.INIT_RAM_08 = 256'hDEC0C0C2687868626878686266666666C0C0C0C2667C6666FEC6C66CDEDEC6C6;
defparam prom_inst_1.INIT_RAM_09 = 256'hC6C6C6C6CEDEFEF6C3DBFFFF6060606078786C660C0C0C0C18181818C6FEC6C6;
defparam prom_inst_1.INIT_RAM_0A = 256'hDBC3C3C3C3C3C3C3C6C6C6C6181818990C3860C66C7C6666C6C6C6C6607C6666;
defparam prom_inst_1.INIT_RAM_0B = 256'h00000000000000000C0C0C0C3870E0C03030303030180C86183C66C318183C66;
defparam prom_inst_1.INIT_RAM_0C = 256'hCCCC760060F06064FEC67C00CC6C3C0CC0C67C00666C78607C0C780000000000;
defparam prom_inst_1.INIT_RAM_0D = 256'hC6C67C006666DC00DBFFE60018181818786C666006060E001818380066766C60;
defparam prom_inst_1.INIT_RAM_0E = 256'hC3C3C300C3C3C300CCCCCC003030FC3060C67C006676DC00CCCC76006666DC00;
defparam prom_inst_1.INIT_RAM_0F = 256'hC66C381000000000180E1818180018181870181818CCFE00C6C6C6003C66C300;

pROM prom_inst_2 (
    .DO(dout[95:64]),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({gw_gnd,gw_gnd,ad[6:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_2.READ_MODE = 1'b0;
defparam prom_inst_2.BIT_WIDTH = 32;
defparam prom_inst_2.RESET_MODE = "SYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'h0000183C3C18187E3C1818E70010387C10387CFE7EFFFFE77E81819900000000;
defparam prom_inst_2.INIT_RAM_01 = 256'h1818DB3CE6E76763E0F0703018187E1878CCCCCCFFC399BD003C6642FFFFE7C3;
defparam prom_inst_2.INIT_RAM_02 = 256'h7E183C7EFEFEFEFEC60C386C1B1B1B1B6666006600183C7E02060E1E80C0E0F0;
defparam prom_inst_2.INIT_RAM_03 = 256'h0010383800FEFE7C000024660000FEC0000030600000180C183C7E1818181818;
defparam prom_inst_2.INIT_RAM_04 = 256'h0000000076CCCCCC86C660307CC686066C6CFE6C000000001818001800000000;
defparam prom_inst_2.INIT_RAM_05 = 256'h80C06030181800000000000018181800000018180000663C30180C0C0C183030;
defparam prom_inst_2.INIT_RAM_06 = 256'h303030307CC6C6C67CC606061E0C0C0C7CC60606FEC6C0607E1818187CC6C6E6;
defparam prom_inst_2.INIT_RAM_07 = 256'h181800186030180C0000007E060C18303018180000181800780C06067CC6C6C6;
defparam prom_inst_2.INIT_RAM_08 = 256'h3A66C6C6F0606060FE666260F86C66663C66C2C0FC666666C6C6C6C67CC0DCDE;
defparam prom_inst_2.INIT_RAM_09 = 256'h7CC6C6C6C6C6C6C6C3C3C3C3FE666260E666666C78CCCCCC3C181818C6C6C6C6;
defparam prom_inst_2.INIT_RAM_0A = 256'h6666FFDB183C66C37CC6C6C63C1818187CC6C606E66666667CDED6C6F0606060;
defparam prom_inst_2.INIT_RAM_0B = 256'h00000000000000003C0C0C0C02060E1C3C303030FFC3C1603C181818C3C3663C;
defparam prom_inst_2.INIT_RAM_0C = 256'h7CCCCCCCF06060607CC6C0C076CCCCCC7CC6C0C07C66666676CCCCCC00000000;
defparam prom_inst_2.INIT_RAM_0D = 256'h7CC6C6C666666666DBDBDBDB3C181818E6666C78060606063C181818E6666666;
defparam prom_inst_2.INIT_RAM_0E = 256'h66FFDBDB183C66C376CCCCCC1C3630307CC60C38F06060607CCCCCCC7C666666;
defparam prom_inst_2.INIT_RAM_0F = 256'h00FEC6C60000000070181818181818180E181818FEC660307EC6C6C6C3663C18;

pROM prom_inst_3 (
    .DO(dout[127:96]),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({gw_gnd,gw_gnd,ad[6:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_3.READ_MODE = 1'b0;
defparam prom_inst_3.BIT_WIDTH = 32;
defparam prom_inst_3.RESET_MODE = "SYNC";
defparam prom_inst_3.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_01 = 256'h00000000000000C0000000000000000000000000FFFFFFFF00000000FFFFFFFF;
defparam prom_inst_3.INIT_RAM_02 = 256'h00000000000000000000007C0000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_04 = 256'h0000000000000000000000000000181800000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_05 = 256'h0000000000000000000000000000003000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_0A = 256'h00000000000000000000000000000000000000000000000000000E0C00000000;
defparam prom_inst_3.INIT_RAM_0B = 256'h0000FF0000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_0C = 256'h0078CC0C00000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000003C66660000000000000000;
defparam prom_inst_3.INIT_RAM_0E = 256'h000000000000000000000000000000000000000000000000001E0C0C00F06060;
defparam prom_inst_3.INIT_RAM_0F = 256'h00000000000000000000000000000000000000000000000000F80C0600000000;

endmodule //Gowin_pROM
